/***********************************************************************
 * A SystemVerilog top-level netlist to connect testbench to DUT
 **********************************************************************/

module top;
  //directiva de compilator - seteaza timpul de simulare (rezolutie, pasul)
  timeunit 1ns/1ns;

  // user-defined types are defined in instr_register_pkg.sv
  import instr_register_pkg::*;

  // clock variables
  logic clk;
  logic test_clk;

  // interconnecting signals
  logic          reset_n;


  tb_ifc tbifc();  // instantiate testbench and connect ports

  instr_register dut(
                    .tbif(tbifc.DUT),
                    .clk (clk), 
                    .reset_n (reset_n));

  instr_register_test test(
                          .tbif(tbifc.TEST),
                          .clk (test_clk), 
                          .reset_n (reset_n));

  // clock oscillators
  initial begin
    clk <= 0;
    forever #5  clk = ~clk;
  end

  initial begin
    test_clk <=0;
    // offset test_clk edges from clk to prevent races between
    // the testbench and the design
    #4 forever begin
      #2ns test_clk = 1'b1;
      #8ns test_clk = 1'b0;
    end
  end

endmodule: top
